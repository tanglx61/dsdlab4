library verilog;
use verilog.vl_types.all;
entity g58_rules_test_vlg_vec_tst is
end g58_rules_test_vlg_vec_tst;
