library verilog;
use verilog.vl_types.all;
entity g58_rules_test_vlg_check_tst is
    port(
        legal_play      : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end g58_rules_test_vlg_check_tst;
